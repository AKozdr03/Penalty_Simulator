/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Authors: Andrzej Kozdrowski, Aron Lampart
 * Description:
 * End screen controler.
 */

 module end_screen(
    input wire clk,
    input wire rst

    );
       
      
endmodule