/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Authors: Andrzej Kozdrowski, Aron Lampart
 * Description:
 * Drawing gloves on the screen.
 */

 module draw_gloves(
    input wire clk,
    input wire rst,
    input wire [11:0] xpos, ypos

);
   
  
endmodule