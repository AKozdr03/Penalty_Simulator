/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Author: Andrzej Kozdrowski
 *
 * Description:
 * 256 characters :).
 */

module char_16x16(
    input wire clk,
    input logic [7:0] char_xy,
    
    output logic [6:0] char_code
);
    logic [6:0] data;

always_ff @(posedge clk)
    char_code <= data;

always_comb begin
    case(char_xy) 
        8'h00: data = "W";
        8'h01: data = "I";
        8'h02: data = "E";
        8'h03: data = "L";
        8'h04: data = "E";
        8'h05: data = " ";  
        8'h06: data = "R";
        8'h07: data = "Z";
        8'h08: data = "E";
        8'h09: data = "C";
        8'h0a: data = "Z";
        8'h0b: data = "Y";
        8'h0c: data = " ";
        8'h0d: data = " ";
        8'h0e: data = " ";
        8'h0f: data = " ";
        8'h10: data = "M";
        8'h11: data = "O";
        8'h12: data = "Z";
        8'h13: data = "E";
        8'h14: data = "M";
        8'h15: data = "Y";
        8'h16: data = " ";
        8'h17: data = " ";
        8'h18: data = " ";
        8'h19: data = " ";
        8'h1a: data = " ";
        8'h1b: data = " ";
        8'h1c: data = " ";
        8'h1d: data = " ";
        8'h1e: data = " ";
        8'h1f: data = " ";
        8'h20: data = "Z";
        8'h21: data = "A";
        8'h22: data = "C";
        8'h23: data = "H";
        8'h24: data = "O";
        8'h25: data = "W";
        8'h26: data = "A";
        8'h27: data = "C";
        8'h28: data = " ";
        8'h29: data = "L";
        8'h2a: data = "U";
        8'h2b: data = "B";
        8'h2c: data = " ";
        8'h2d: data = " ";
        8'h2e: data = " ";
        8'h2f: data = " ";

        8'h30: data = "Z";
        8'h31: data = "N";
        8'h32: data = "I";
        8'h33: data = "S";
        8'h34: data = "Z";
        8'h35: data = "C";  
        8'h36: data = "Z";
        8'h37: data = "Y";
        8'h38: data = "C";
        8'h39: data = " ";
        8'h3a: data = "J";
        8'h3b: data = "E";
        8'h3c: data = "D";
        8'h3d: data = "N";
        8'h3e: data = "Y";
        8'h3f: data = "M";
        8'h40: data = "Z";
        8'h41: data = " ";
        8'h42: data = "P";
        8'h43: data = "O";
        8'h44: data = "Z";
        8'h45: data = "O";
        8'h46: data = "R";
        8'h47: data = "U";
        8'h48: data = " ";
        8'h49: data = " ";
        8'h4a: data = " ";
        8'h4b: data = " ";
        8'h4c: data = " ";
        8'h4d: data = " ";
        8'h4e: data = " ";
        8'h4f: data = " ";
        8'h50: data = "N";
        8'h51: data = "I";
        8'h52: data = "E";
        8'h53: data = "W";
        8'h54: data = "A";
        8'h55: data = "Z";
        8'h56: data = "N";
        8'h57: data = "Y";
        8'h58: data = "M";
        8'h59: data = " ";
        8'h5a: data = "G";
        8'h5b: data = "E";
        8'h5c: data = "S";
        8'h5d: data = "T";
        8'h5e: data = "E";
        8'h5f: data = "M";        

        8'h60: data = "~";
        8'h61: data = "P";
        8'h62: data = "A";
        8'h63: data = "U";
        8'h64: data = "L";
        8'h65: data = "0";  
        8'h66: data = " ";
        8'h67: data = "C";
        8'h68: data = "O";
        8'h69: data = "E";
        8'h6a: data = "L";
        8'h6b: data = "H";
        8'h6c: data = "O";
        8'h6d: data = " ";
        8'h6e: data = " ";
        8'h6f: data = " ";
        8'h70: data = " ";
        8'h71: data = " ";
        8'h72: data = " ";
        8'h73: data = " ";
        8'h75: data = " ";
        8'h76: data = " ";
        8'h77: data = " ";
        8'h78: data = " ";
        8'h79: data = " ";
        8'h7a: data = " ";
        8'h7b: data = " ";
        8'h7c: data = " ";
        8'h7d: data = " ";
        8'h7e: data = " ";
        8'h7f: data = " ";
        8'h80: data = " ";
        8'h81: data = " ";
        8'h82: data = " ";
        8'h83: data = " ";
        8'h84: data = " ";
        8'h85: data = " ";
        8'h86: data = " ";
        8'h87: data = " ";
        8'h88: data = " ";
        8'h89: data = " ";
        8'h8a: data = " ";
        8'h8b: data = " ";
        8'h8c: data = " ";
        8'h8d: data = " ";
        8'h8e: data = " ";
        8'h8f: data = " ";
        
        8'h90: data = " ";
        8'h91: data = " ";
        8'h92: data = " ";
        8'h93: data = " ";
        8'h94: data = " ";
        8'h95: data = " ";  
        8'h96: data = " ";
        8'h97: data = " ";
        8'h98: data = " ";
        8'h99: data = " ";
        8'h9a: data = " ";
        8'h9b: data = " ";
        8'h9c: data = " ";
        8'h9d: data = " ";
        8'h9e: data = " ";
        8'h9f: data = " ";
        8'ha0: data = " ";
        8'ha1: data = " ";
        8'ha2: data = " ";
        8'ha3: data = " ";
        8'ha5: data = " ";
        8'ha6: data = " ";
        8'ha7: data = " ";
        8'ha8: data = " ";
        8'ha9: data = " ";
        8'haa: data = " ";
        8'hab: data = " ";
        8'hac: data = " ";
        8'had: data = " ";
        8'hae: data = " ";
        8'haf: data = " ";
        8'hb0: data = " ";
        8'hb1: data = " ";
        8'hb2: data = " ";
        8'hb3: data = " ";
        8'hb4: data = " ";
        8'hb5: data = " ";
        8'hb6: data = " ";
        8'hb7: data = " ";
        8'hb8: data = " ";
        8'hb9: data = " ";
        8'hba: data = " ";
        8'hbb: data = " ";
        8'hbc: data = " ";
        8'hbd: data = " ";
        8'hbe: data = " ";
        8'hbf: data = " ";
        8'hc0: data = " ";
        8'hc1: data = " ";
        8'hc2: data = " ";
        8'hc3: data = " ";
        8'hc4: data = " ";
        8'hc5: data = " ";  
        8'hc6: data = " ";
        8'hc7: data = " ";
        8'hc8: data = " ";
        8'hc9: data = " ";
        8'hca: data = " ";
        8'hcb: data = " ";
        8'hcc: data = " ";
        8'hcd: data = " ";
        8'hce: data = " ";
        8'hcf: data = " ";
        8'hd0: data = "P";
        8'hd1: data = "O";
        8'hd2: data = "Z";
        8'hd3: data = "D";
        8'hd4: data = "R";
        8'hd5: data = "A";
        8'hd6: data = "W";
        8'hd7: data = "I";
        8'hd8: data = "A";
        8'hd9: data = "M";
        8'hda: data = " ";
        8'hdb: data = " ";
        8'hdc: data = " ";
        8'hdd: data = " ";
        8'hde: data = " ";
        8'hdf: data = " ";
        8'he0: data = "A";
        8'he1: data = "N";
        8'he2: data = "D";
        8'he3: data = "R";
        8'he4: data = "Z";
        8'he5: data = "E";
        8'he6: data = "J";
        8'he7: data = " ";
        8'he8: data = " ";
        8'he9: data = " ";
        8'hea: data = " ";
        8'heb: data = " ";
        8'hec: data = " ";
        8'hed: data = " ";
        8'hee: data = " ";
        8'hef: data = " ";       
        8'hf0: data = "K";
        8'hf1: data = "O";
        8'hf2: data = "Z";
        8'hf3: data = "D";
        8'hf4: data = "R";
        8'hf5: data = "O";
        8'hf6: data = "W";
        8'hf7: data = "S";
        8'hf8: data = "K";
        8'hf9: data = "I";
        8'hfa: data = " ";
        8'hfb: data = " ";
        8'hfc: data = " ";
        8'hfd: data = " ";
        8'hfe: data = " ";
        8'hff: data = " ";   
    endcase
        end

endmodule