/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Authors: Andrzej Kozdrowski, Aron Lampart
 * Description:
 * Shooter screen controler.
 */

 module shooter_screen(
    input wire clk,
    input wire rst
);
   
  
endmodule