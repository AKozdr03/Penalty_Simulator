/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Authors: Andrzej Kozdrowski, Aron Lampart
 * Description:
 * Drawing keeper on the screen.
 */

 module draw_keeper(
    input wire clk,
    input wire rst
);
   
  
endmodule