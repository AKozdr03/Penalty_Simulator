/**
 * Copyright (C) 2024  AGH University of Science and Technology
 * MTM UEC2
 * Authors: Andrzej Kozdrowski, Aron Lampart
 * Description:
 * Ball controller.
 */

 module ball_control(
    input wire clk, rst
);



endmodule